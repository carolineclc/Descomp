library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity ExtensorSinal IS
   port ( 

          Dado_in  : in std_logic_vector(15 downto 0);
          Dado_out : out std_logic_vector(31 downto 0)

        );
end entity;

architecture assincrona OF ExtensorSinal IS
signal extensao : std_logic_vector(15 downto 0); 

begin
	
	extensao <= (others => Dado_in(15));

  Dado_out <= extensao & Dado_in ;

end architecture;