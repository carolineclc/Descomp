library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
        tmp(0)  := "1001000001110";   -- Desta posicao para baixo, é necessário acertar os valores
        tmp(1)  := "0110000000101";	  -- 
        tmp(2)  := "0111000001001";
        tmp(3)  := "0000000000000";
        tmp(4)  := "0000000000000";
        tmp(5)  := "0100000000101";
        tmp(6)  := "0101100000000";
		  tmp(7)  := "1000100000000";
		  tmp(8)  := "0110000000010";
		  tmp(9)  := "0000000000000";
		  tmp(10) := "0100000000100";
		  tmp(11) := "1000100000000";
		  tmp(12) := "0111000000011";
		  tmp(13) := "0110000001101";
		  tmp(14) := "0000000000000";
		  tmp(15) := "1010000000000";
      
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;