library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  
  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
		  


  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := x"4" & '0' & x"00";	-- LDI $0
tmp(1) := x"5" & '1' & x"20";	-- STA @288
tmp(2) := x"5" & '1' & x"21";	-- STA @289
tmp(3) := x"5" & '1' & x"22";	-- STA @290
tmp(4) := x"5" & '1' & x"23";	-- STA @291
tmp(5) := x"5" & '1' & x"24";	-- STA @292
tmp(6) := x"5" & '1' & x"25";	-- STA @293
tmp(7) := x"5" & '1' & x"00";	-- STA @256
tmp(8) := x"5" & '1' & x"01";	-- STA @257
tmp(9) := x"5" & '1' & x"02";	-- STA @258
tmp(10) := x"5" & '1' & x"FF";	-- STA @511 	#LIMPA FLAG DO BOTAO KEY0
tmp(11) := x"5" & '1' & x"FE";	-- STA @510 	#LIMPA FLAG DO BOTAO KEY1
tmp(12) := x"5" & '0' & x"00";	-- STA @0 	#ARMAZENA O VALOR DO ACUMULADOR EM MEM[0] (UNIDADES)
tmp(13) := x"5" & '0' & x"01";	-- STA @1 	#ARMAZRNA O VALOR DO ACUMULADOR EM MEM [1] (DEZENAS)
tmp(14) := x"5" & '0' & x"02";	-- STA @2 	#ARMAZENA O VALOR DO ACUMULADOR EM MEM [2] (CENENAS)
tmp(15) := x"5" & '0' & x"05";	-- STA @5 	#ARMAZENA O VALOR DO ACUMULADOR EM MEM [5] (FLAG UNIDADE)
tmp(16) := x"5" & '0' & x"06";	-- STA @6 	#ARMAZENA O VALOR DO ACUMULADOR EM MEM [6] (LIMITE)
tmp(17) := x"5" & '0' & x"07";	-- STA @7 	#ARMAZENA O VALOR DO ACUMULADOR EM MEM [7] (FLAG LIMITE)
tmp(18) := x"5" & '0' & x"03";	-- STA @3 	# CONSTANTE 0
tmp(19) := x"4" & '0' & x"01";	-- LDI $1
tmp(20) := x"5" & '0' & x"04";	-- STA @4 	#CONSTANTE 1
tmp(21) := x"1" & '1' & x"61";	-- LDA @353 	#LE O VALOR DO BOTAO DE  KEY0
tmp(22) := x"8" & '0' & x"03";	-- CEQ @3 	#COMPARA SE O VALOR DE KEY0 IGUAL A 0
tmp(23) := x"7" & '0' & x"19";	-- JEQ @cont 	#SE KEY0 NAO FOI PRESSIONADO CONTUNA NO LACO
tmp(24) := x"9" & '0' & x"28";	-- JSR @incremento 	#SE KEY0 FOI PRESSIONADO ENTRA NA SUBROTINA DE INREMENTO
tmp(25) := x"9" & '0' & x"33";	-- JSR @ display
tmp(26) := x"1" & '1' & x"60";	-- LDA @352 	#LE O VALOR DO BOTAO DE  KEY1
tmp(27) := x"8" & '0' & x"03";	-- CEQ @3 	#COMPARA SE O VALOR DE KEY0 IGUAL A 0
tmp(28) := x"7" & '0' & x"19";	-- JEQ @cont 	#SE KEY1 NAO FOI PRESSIONADO VOLTA PARA O INICIO
tmp(29) := x"9" & '0' & x"2E";	-- JSR @limite 	#SE KEY0 FOI PRESSIONADO ENTRA NA SUBROTINA DE INREMENTO
tmp(30) := x"1" & '0' & x"06";	-- LDA @6 	#PEGA VALOR DE LIMITE
tmp(31) := x"5" & '1' & x"22";	-- STA @290 	#DISPLAY VALOR DE LIMITE EM HEX2
tmp(32) := x"1" & '0' & x"00";	-- LDA @0 	#PEGA O VALOR DAS UNIDADES
tmp(33) := x"8" & '0' & x"06";	-- CEQ @6 	#COMPARA COM O VALOR DO LIMITE
tmp(34) := x"7" & '0' & x"36";	-- JEQ @final 	#SE FOR IGUAL VAI NO FINAL
tmp(35) := x"1" & '1' & x"64";	-- LDA @356 	#PEGA O VALOR DO BOTAO FPGA RESET
tmp(36) := x"8" & '0' & x"03";	-- CEQ @3 	#COMPARA SE O VALOR DE FPGA RESET FOI PRESSIONADO
tmp(37) := x"7" & '0' & x"27";	-- JEQ @cont3 	#SE O BOTAO NAO FOI PRESSIONADO CONTINUA NO LACO
tmp(38) := x"9" & '0' & x"00";	-- JSR @limpeza 	#SE O BOTAO FOI PRESSIONADO ELE FAZ A LIMPEZA DAS VARIAVEIS
tmp(39) := x"6" & '0' & x"15";	-- JMP @inicio
tmp(40) := x"1" & '0' & x"03";	-- LDA @3
tmp(41) := x"5" & '1' & x"FE";	-- STA @510 	#LIMPA A FLAG DO BOTAO KEY0
tmp(42) := x"1" & '0' & x"04";	-- LDA @4 	#ARMAZENA A CONSTANTE NO REGISTRADOR
tmp(43) := x"2" & '0' & x"00";	-- SOMA @0 	#SOMA A CONSTANTE NO VALOR DAS UNIDADES
tmp(44) := x"5" & '0' & x"00";	-- STA @0 	#ARMAZENA O NOVO VALOR NAS UNIDADES
tmp(45) := x"A" & '0' & x"00";	-- RET
tmp(46) := x"1" & '1' & x"40";	-- LDA @320 	#PEGA OS VALORES DA CHAVE
tmp(47) := x"5" & '0' & x"06";	-- STA @6 	#ARMAZENA NA VARIAVEL DE MEM[6]
tmp(48) := x"4" & '0' & x"01";	-- LDI $1 	#CONSTANTE 1
tmp(49) := x"5" & '1' & x"01";	-- STA @257 	#ACENDE LED8 INDICANDO QUE LIMITE FOI DEFINIDO
tmp(50) := x"A" & '0' & x"00";	-- RET
tmp(51) := x"1" & '0' & x"00";	-- LDA @0 	#PEGA O VALOR DAS UNIDADES
tmp(52) := x"5" & '1' & x"20";	-- STA @288 	#ESCREVE O VALOR NO DISPLAY HEX0
tmp(53) := x"A" & '0' & x"00";	-- RET
tmp(54) := x"4" & '0' & x"01";	-- LDI $1
tmp(55) := x"5" & '1' & x"02";	-- STA @258 	#ACENDE LED9 INDICANDO QUE LIMITE FOI ATINGIDO
tmp(56) := x"6" & '0' & x"15";	-- JMP @inicio





        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;